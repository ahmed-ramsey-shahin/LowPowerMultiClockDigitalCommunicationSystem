module GrayCodeEncoder (
    input  wire [4:0] x,
    output reg  [4:0] y
);
    always @(*) begin
        case (x)
            5'd0:  y = 5'b00000;
            5'd1:  y = 5'b00001;
            5'd2:  y = 5'b00011;
            5'd3:  y = 5'b00010;
            5'd4:  y = 5'b00110;
            5'd5:  y = 5'b00111;
            5'd6:  y = 5'b00101;
            5'd7:  y = 5'b00100;
            5'd8:  y = 5'b01100;
            5'd9:  y = 5'b01101;
            5'd10: y = 5'b01111;
            5'd11: y = 5'b01110;
            5'd12: y = 5'b01010;
            5'd13: y = 5'b01011;
            5'd14: y = 5'b01001;
            5'd15: y = 5'b01000;
            5'd16: y = 5'b11000;
            5'd17: y = 5'b11001;
            5'd18: y = 5'b11011;
            5'd19: y = 5'b11010;
            5'd20: y = 5'b11110;
            5'd21: y = 5'b11111;
            5'd22: y = 5'b11101;
            5'd23: y = 5'b11100;
            5'd24: y = 5'b10100;
            5'd25: y = 5'b10101;
            5'd26: y = 5'b10111;
            5'd27: y = 5'b10110;
            5'd28: y = 5'b10010;
            5'd29: y = 5'b10011;
            5'd30: y = 5'b10001;
            5'd31: y = 5'b10000;
        endcase
    end
endmodule
